`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AIST
// Engineer: Junichi Sakamoto
// 
// Create Date: 2024/12/12
// Module Name: tb_ML_KEM.sv
// Tool Versions: Vivado 2024.1
//////////////////////////////////////////////////////////////////////////////////



module tb_ML_KEM;
    localparam integer
        CYCLE = 10,
        DELAY = 1,
        N_LOOP = 20;

    import TYPES_KEM::*;

    reg clk_i, rst_n_i, run_i;
    kem_mode_t mode_i;

    always begin
        #(CYCLE/2) clk_i <= ~clk_i;
    end

    ML_KEM dut (
        .clk_i,
        .rst_n_i,
        .run_i,
        .mode_i
    );

    /*-------------------------------------------
    Test
    -------------------------------------------*/
    initial begin
        clk_i <= 1;
        rst_n_i <= 1;
        #DELAY;
        #100
        rst_n_i <= 0;
        run_i <= 0;
        mode_i <='0;
        #100
        rst_n_i <= 1;
        #100;
        mode_i <= 3'b100;
        run_i <= 1;
        #CYCLE;
        run_i <= 0;

        #1000; 
        //$finish;
    end

endmodule


/*
TV
d = b54b1dbadaba7e84d22ec86169e8702609b165097a072e3b0d1d2fca08409c84
rho = 44359356139e288ce59d819df1b344621e13f705942edf2b8c144eda3eb6846e (little endian)
sigma = 8568575ebf9c1b52642964f3aea51aa87ae9f55a60106713ada487f71a6d5398 (little endian)

A
['0xaab', '0x8b5', '0xb49', '0x7d3', '0x37a', '0x5a5', '0x2d9', '0x83f', '0xb73', '0x22b', '0xcdc', '0x1f6', '0x51', '0x555', '0x8f9', '0xb9d', '0xc2f', '0xabf', '0xbb7', '0xbb6', '0x260', '0xaa2', '0xba6', '0xa2d', '0x120', '0xc06', '0x7de', '0x4b0', '0x757', '0xcb6', '0x3b8', '0xc12', '0x6b3', '0xb27', '0x866', '0x5e2', '0x956', '0x94c', '0x6', '0x39a', '0x900', '0xc19', '0x3cb', '0x872', '0x33a', '0x563', '0x305', '0x97', '0x752', '0xbf4', '0x4d3', '0x42', '0xcb3', '0xb87', '0x3f2', '0x110', '0x251', '0xb44', '0x569', '0xc4e', '0x66d', '0x309', '0x743', '0x31c', '0xc95', '0x9ec', '0x81f', '0x586', '0x7a6', '0x92c', '0x3a', '0x7db', '0xc18', '0x63e', '0xae0', '0xbd0', '0x73', '0x4e1', '0x1a6', '0x53a', '0xb5', '0x6fe', '0x7d3', '0x1a1', '0x252', '0x1ca', '0x369', '0xb', '0x7f1', '0x4c1', '0xca4', '0x588', '0x2c4', '0xb68', '0x440', '0x898', '0x245', '0x77', '0x59d', '0x6e7', '0xb', '0x588', '0x66f', '0x323', '0x91a', '0xc33', '0x3b5', '0x2a5', '0xb09', '0x3ab', '0x2de', '0x333', '0xb11', '0x887', '0x5ff', '0xb65', '0x143', '0x7b7', '0xac0', '0xe1', '0x9ee', '0xa29', '0x9d5', '0xa9d', '0xb26', '0x4a9', '0x2db', '0x115', '0x14a', '0xb3a', '0x3aa', '0xb7b', '0x42a', '0xbf6', '0x2ee', '0x19e', '0x75c', '0x4b9', '0x6a8', '0xa6e', '0x16f', '0x118', '0xe1', '0x4bc', '0x4d0', '0x9', '0x8d4', '0x8e6', '0x13d', '0x202', '0x211', '0x1f2', '0x264', '0x4f0', '0x7d5', '0xcb0', '0x455', '0xb50', '0xc0c', '0x93d', '0x687', '0xa1f', '0x6b3', '0xbe8', '0x807', '0x3ca', '0x51a', '0x36c', '0x81a', '0x368', '0x6a9', '0x716', '0x3d9', '0x924', '0x31d', '0x3f4', '0x163', '0x54d', '0xc2b', '0x28d', '0x416', '0x83d', '0xbf5', '0x200', '0xbb', '0x511', '0x72c', '0xc28', '0xc5f', '0xc99', '0xa88', '0x129', '0x61e', '0x791', '0xb04', '0xbab', '0x272', '0x9d0', '0x529', '0xa65', '0x313', '0x841', '0x97e', '0x51a', '0x841', '0xb7f', '0x18', '0xce7', '0x73c', '0x33a', '0x79', '0xbcc', '0xa69', '0xbf6', '0x391', '0x43a', '0x378', '0x333', '0xcf2', '0x528', '0x473', '0xcfb', '0x998', '0x1c4', '0x7d', '0x734', '0x5fd', '0xbf4', '0xa1e', '0x9ce', '0x64b', '0x261', '0x1b6', '0x481', '0x71f', '0x84d', '0xa5c', '0x43b', '0xce1', '0x260', '0xb7c', '0xabc', '0x4dd', '0xc7', '0x740', '0x373', '0x442', '0x267', '0x1b0', '0x203', '0x587', '0x567', '0x55a', '0x67f', '0x188', '0x961']
['0x930', '0x44a', '0x445', '0x89c', '0x268', '0x96a', '0x39b', '0x6c3', '0xc96', '0x6ef', '0x5d4', '0xc53', '0x292', '0x709', '0x4eb', '0x49', '0xcf8', '0xa59', '0xb9f', '0xbb1', '0xc6e', '0xa9d', '0x3b7', '0x72a', '0x822', '0x1b9', '0xb50', '0xaf8', '0xe6', '0x1a5', '0x5f0', '0xa73', '0xa18', '0xce7', '0xb0b', '0x2c1', '0x173', '0xa81', '0xa1a', '0x4e6', '0xbc9', '0x5c4', '0x78', '0xbbb', '0x768', '0xc81', '0x2c2', '0x442', '0x4a8', '0x55c', '0x1ac', '0x306', '0x381', '0x279', '0x369', '0x97c', '0xa52', '0x268', '0x859', '0x33f', '0x77f', '0x95c', '0xb6d', '0x643', '0xf', '0x82c', '0x581', '0x144', '0xa0a', '0x15e', '0x4f4', '0xa3e', '0x107', '0xa12', '0x6bf', '0x6f0', '0x7b8', '0x314', '0x943', '0x611', '0x4e4', '0x4ff', '0xbe1', '0x29c', '0xad4', '0x123', '0x2e7', '0x311', '0x478', '0x219', '0x99a', '0xce3', '0xc1e', '0x1bd', '0x759', '0x264', '0x957', '0xb6c', '0x320', '0x63f', '0x9cb', '0xb4a', '0x2ca', '0xc25', '0x658', '0xc0c', '0x43f', '0xccf', '0x765', '0x2e7', '0x56b', '0xb31', '0x28a', '0x393', '0x549', '0x35', '0x3ad', '0x77d', '0xcef', '0xc99', '0x248', '0x8fd', '0xcd0', '0xaa8', '0xb77', '0x779', '0x161', '0x2b0', '0x31', '0x8b6', '0x556', '0x601', '0xc30', '0xad9', '0x528', '0x7e4', '0xb26', '0x697', '0x6fb', '0x828', '0x454', '0x89e', '0x317', '0x85c', '0xc1b', '0x8fd', '0x9c4', '0x306', '0x934', '0x20', '0x568', '0x47', '0x733', '0x4be', '0x6cc', '0xf1', '0x98b', '0xc8a', '0xad4', '0x915', '0xa38', '0x200', '0xa3f', '0x62a', '0xbbe', '0x8c7', '0xbcf', '0x3a8', '0x5f4', '0x11', '0x32e', '0x54a', '0xc59', '0x4a1', '0x36e', '0x739', '0x7fd', '0x670', '0x5a2', '0x357', '0xe7', '0x704', '0xaa0', '0x40c', '0xd9', '0x97c', '0x473', '0xadb', '0x782', '0xb99', '0x527', '0x58', '0xadf', '0x5a6', '0x365', '0x318', '0xa6f', '0x84', '0x8cc', '0x423', '0x64b', '0x581', '0x794', '0x3a', '0xb98', '0xa7d', '0x85', '0xbe6', '0x7f', '0x693', '0x25d', '0x19a', '0x6e7', '0xb7b', '0x134', '0x3d0', '0x900', '0x627', '0x34c', '0x2bb', '0x314', '0x905', '0xa12', '0x2f8', '0x9dd', '0xc71', '0x3ba', '0x78d', '0x21a', '0x8bf', '0x9a4', '0x547', '0xb1a', '0x322', '0x8d3', '0xb11', '0x9d1', '0x5c1', '0x480', '0x2bb', '0x87f', '0x9ea', '0x5f3', '0x99f', '0xcf6', '0xbaf', '0x1c0', '0x2ed', '0x669', '0x839', '0xc74', '0x4bc', '0x5eb', '0x15d', '0x5df', '0x82b']
['0x494', '0x2ff', '0x872', '0xc8e', '0x22b', '0x4c5', '0x522', '0xc3', '0x8c2', '0x56d', '0x616', '0x654', '0xc26', '0x1df', '0x817', '0xb70', '0x779', '0x6bc', '0x8a0', '0x134', '0xb4', '0xb1e', '0x72f', '0x4da', '0x885', '0x845', '0xbb7', '0x40a', '0x55d', '0x7bf', '0x9f2', '0x536', '0x3ea', '0x407', '0x650', '0x5ce', '0x5a3', '0x851', '0x88a', '0x308', '0xa2c', '0x12d', '0x6fa', '0x4b3', '0x196', '0x1c5', '0x12c', '0x1ce', '0x469', '0x7c2', '0xac5', '0x89', '0x8c3', '0x405', '0xc75', '0x7fe', '0xc76', '0x2cb', '0x3d3', '0x922', '0x17b', '0x15', '0x824', '0x691', '0x3f8', '0x230', '0x7f3', '0x95a', '0x668', '0x1e', '0x6ef', '0xc75', '0x5f2', '0x6b7', '0x61d', '0x310', '0x18b', '0x1c7', '0x1d4', '0x920', '0xbc7', '0x11', '0x788', '0x4b0', '0xa11', '0x9b7', '0x82', '0x99b', '0x18a', '0x6ba', '0xef', '0x85e', '0x482', '0xcf8', '0x1d0', '0x90d', '0xa03', '0x5ca', '0x613', '0x6fd', '0x31d', '0x363', '0x971', '0x1bf', '0x5ef', '0x6de', '0xc04', '0x42f', '0x8d5', '0x602', '0x9ac', '0xc28', '0x308', '0x2f6', '0x8aa', '0x892', '0x521', '0xa3e', '0xb81', '0x72a', '0x1b1', '0x4fb', '0x6f5', '0xcb9', '0x8c7', '0x967', '0x395', '0xa1b', '0xb61', '0x64b', '0x541', '0x157', '0xc2', '0x54', '0x342', '0xa7f', '0x8c2', '0x207', '0xa3b', '0x9de', '0x901', '0x4dc', '0xa8', '0x9dc', '0xc42', '0x1e0', '0xb22', '0x62a', '0x698', '0x64', '0x2cd', '0x1e8', '0x5ab', '0x40c', '0x376', '0x83b', '0x998', '0x957', '0x143', '0x47c', '0x9ab', '0xc92', '0x39e', '0x280', '0x8db', '0x908', '0x93c', '0xc89', '0x7cd', '0x78e', '0x3ee', '0x984', '0xb8b', '0xc28', '0xc06', '0x721', '0xb9', '0xc75', '0x102', '0x90c', '0xf2', '0xb80', '0x10c', '0x500', '0xaab', '0xb6c', '0x51b', '0xa91', '0x176', '0x6e6', '0x135', '0xc7b', '0x6e0', '0xf0', '0x2fc', '0x9ad', '0x453', '0x992', '0xbc', '0x1f6', '0x4ed', '0x839', '0x77', '0x37d', '0x1bf', '0x18f', '0x7ef', '0x8c2', '0x233', '0x10', '0x7d1', '0xca0', '0x2b9', '0xa23', '0x91a', '0xc57', '0xa0', '0x137', '0x16a', '0x723', '0x933', '0x2f0', '0x4b', '0x4c7', '0x139', '0xc84', '0x339', '0x4f', '0x24f', '0x8a', '0xe5', '0x401', '0x7ef', '0x71', '0x1e3', '0x685', '0x101', '0x1b0', '0x392', '0x76a', '0x98', '0x11f', '0x899', '0xb1e', '0x806', '0x8', '0x60d', '0x403', '0x394', '0x516', '0x84f', '0x6de', '0x844', '0xb00', '0x745', '0xb']
['0xab', '0x514', '0x1af', '0xa4f', '0x9dd', '0x480', '0x896', '0x7e1', '0x40b', '0x397', '0xba7', '0x401', '0x5e9', '0xc17', '0x40f', '0x341', '0x241', '0xc2b', '0x3f0', '0x862', '0x450', '0xaf4', '0x19c', '0x546', '0xaae', '0x785', '0xbe6', '0x24e', '0x938', '0xc53', '0xa4a', '0x90a', '0x1a6', '0xa80', '0x3e2', '0x260', '0x9d2', '0xc61', '0x8e9', '0xa86', '0x1f4', '0x6b3', '0x254', '0x964', '0x9e4', '0x98a', '0x50d', '0xcc5', '0x3ed', '0x875', '0xc40', '0xb0a', '0x53', '0xc6b', '0xcc8', '0x9e1', '0xc15', '0x4ea', '0xa03', '0x639', '0x800', '0x3bd', '0xa7', '0xa19', '0xd1', '0xcf7', '0x58e', '0xa3', '0x908', '0xb97', '0x943', '0xb66', '0xbb7', '0xaab', '0xbff', '0x732', '0x56d', '0x704', '0x27c', '0xc92', '0xc00', '0x3f6', '0x41d', '0x61c', '0x533', '0xbe7', '0x9c2', '0x304', '0xc41', '0x876', '0x256', '0x507', '0x142', '0x2d5', '0x744', '0x336', '0xce1', '0xb1b', '0xd8', '0x7d6', '0x945', '0xbf6', '0xbbc', '0x8b9', '0x1e6', '0x6b8', '0x23b', '0x8d3', '0xc26', '0xae3', '0x33a', '0x65f', '0x521', '0x67f', '0x227', '0xf2', '0xbcc', '0x482', '0x9d7', '0x2f4', '0x5fa', '0xf6', '0x1b2', '0xbce', '0xa57', '0x948', '0xcaa', '0x214', '0x944', '0x8d', '0xc48', '0x58c', '0x2ed', '0xba4', '0x359', '0x4da', '0x667', '0x3eb', '0xc0f', '0x46d', '0x96e', '0x7cf', '0xc89', '0xc31', '0x6f4', '0x10f', '0x784', '0x149', '0x153', '0x8f8', '0x93d', '0x45d', '0x3b7', '0x568', '0x588', '0x75c', '0x6f1', '0x8de', '0x76c', '0x29e', '0x5d1', '0x3', '0xba6', '0x961', '0x76f', '0x251', '0x170', '0xb6f', '0x51b', '0x25', '0x16b', '0xcb9', '0xbad', '0x364', '0x8b7', '0xc81', '0x1cd', '0x177', '0x214', '0xb2f', '0x684', '0xbc7', '0x74b', '0xfa', '0xa99', '0x8d8', '0xb36', '0x6a', '0x390', '0xcb7', '0x362', '0xadd', '0xad5', '0x5a0', '0xcdb', '0xa84', '0xc1f', '0x306', '0x9a3', '0x346', '0x4a7', '0x60', '0x3d7', '0xb8f', '0x6da', '0x4e7', '0xb5b', '0x2a7', '0x9b9', '0x8c9', '0x713', '0xc76', '0xa69', '0x374', '0x5f5', '0x48', '0x79f', '0x6cf', '0xa1', '0xb93', '0x10a', '0x46e', '0x881', '0x616', '0x8ad', '0xd2', '0x190', '0xb0e', '0x4a', '0x5ab', '0xabe', '0x80e', '0xb28', '0xaf', '0xa47', '0x206', '0x67e', '0xa3a', '0x15e', '0x545', '0x902', '0xcd9', '0x724', '0x7d3', '0x4b9', '0xb7d', '0xb7c', '0x47a', '0x35', '0x87d', '0xaf5', '0x6a4', '0x278', '0x9b1', '0x5ac', '0x2bd']

s
['-0x1', '0x1', '0x0', '0x1', '0x1', '0x2', '0x1', '0x1', '-0x1', '-0x1', '-0x1', '0x1', '0x0', '0x0', '-0x1', '-0x2', '0x1', '0x2', '-0x2', '0x1', '0x0', '0x1', '0x0', '0x0', '0x0', '0x1', '0x0', '0x0', '-0x2', '0x1', '0x3', '0x0', '0x1', '0x1', '0x1', '0x1', '-0x1', '-0x2', '-0x1', '-0x1', '0x0', '0x1', '-0x1', '0x1', '-0x2', '0x2', '0x2', '0x1', '-0x1', '0x0', '0x1', '0x2', '0x3', '0x0', '0x1', '-0x2', '0x1', '0x0', '0x1', '0x0', '0x1', '0x0', '0x0', '0x0', '-0x1', '-0x1', '-0x1', '0x0', '-0x1', '-0x1', '-0x1', '-0x2', '0x0', '0x0', '0x1', '-0x1', '-0x1', '0x0', '0x0', '0x1', '0x0', '-0x2', '0x0', '-0x2', '-0x2', '0x0', '0x1', '-0x1', '0x0', '0x1', '0x0', '0x0', '-0x1', '-0x1', '0x1', '0x0', '-0x1', '0x1', '0x1', '0x0', '-0x1', '0x0', '-0x2', '0x0', '-0x2', '-0x1', '-0x2', '-0x1', '0x0', '0x2', '0x1', '0x0', '0x1', '0x2', '-0x1', '0x1', '0x0', '0x2', '-0x1', '0x0', '-0x1', '0x2', '-0x1', '0x1', '0x1', '0x0', '-0x1', '0x0', '-0x1', '0x1', '-0x2', '0x0', '-0x1', '0x0', '0x1', '-0x1', '0x0', '0x1', '0x1', '0x1', '0x0', '0x1', '0x1', '-0x1', '0x1', '0x0', '0x0', '0x2', '-0x2', '-0x1', '0x0', '-0x1', '0x2', '0x0', '0x0', '0x1', '0x1', '0x1', '0x0', '0x2', '0x1', '0x0', '-0x1', '0x1', '0x0', '-0x2', '-0x1', '0x0', '-0x1', '0x1', '0x0', '-0x1', '-0x1', '-0x1', '0x0', '-0x1', '0x0', '0x1', '0x0', '0x0', '-0x3', '-0x1', '0x1', '0x0', '-0x1', '-0x1', '0x0', '0x1', '-0x2', '0x1', '0x1', '-0x1', '0x0', '-0x1', '0x0', '0x2', '0x2', '-0x1', '-0x1', '-0x1', '-0x1', '-0x1', '-0x2', '-0x3', '-0x1', '0x0', '-0x1', '0x0', '0x0', '0x0', '-0x3', '0x0', '0x0', '-0x2', '0x0', '0x2', '0x2', '-0x1', '0x2', '0x0', '-0x1', '0x1', '-0x1', '0x0', '-0x1', '0x1', '-0x2', '0x1', '-0x1', '-0x1', '0x0', '0x0', '-0x1', '-0x1', '0x1', '0x0', '-0x1', '0x0', '0x0', '0x3', '-0x1', '0x0', '-0x1', '0x2', '0x0', '-0x2', '-0x1', '0x0', '0x0', '-0x1', '0x3', '-0x2', '-0x2', '0x0', '0x0', '-0x1']
['-0x2', '0x0', '0x0', '0x0', '0x0', '0x0', '-0x1', '-0x1', '-0x1', '0x1', '-0x1', '-0x1', '-0x1', '-0x1', '0x0', '-0x1', '-0x1', '-0x1', '-0x1', '0x1', '0x2', '0x1', '-0x2', '0x1', '0x1', '-0x1', '0x2', '-0x1', '0x1', '0x0', '0x1', '0x1', '-0x2', '0x1', '-0x1', '0x3', '0x1', '0x1', '0x0', '0x0', '0x0', '0x0', '0x0', '0x0', '0x1', '-0x1', '0x1', '0x1', '0x2', '-0x1', '0x1', '-0x1', '0x1', '0x0', '0x0', '0x1', '0x0', '-0x2', '-0x2', '0x0', '0x2', '0x0', '0x0', '0x0', '0x1', '-0x1', '0x0', '0x0', '-0x1', '0x0', '-0x2', '0x1', '0x2', '-0x1', '0x0', '-0x1', '-0x1', '-0x1', '0x0', '-0x2', '-0x1', '0x1', '-0x2', '0x1', '0x0', '0x3', '-0x1', '-0x1', '0x0', '-0x1', '0x0', '0x0', '-0x1', '0x0', '0x0', '0x0', '0x0', '0x2', '0x0', '0x0', '-0x1', '0x1', '-0x1', '-0x2', '0x0', '0x1', '-0x1', '-0x2', '0x0', '0x0', '0x1', '0x0', '0x0', '-0x2', '-0x1', '0x2', '0x1', '0x1', '-0x2', '0x0', '-0x1', '0x0', '-0x1', '0x1', '-0x1', '0x1', '-0x2', '0x1', '0x0', '-0x2', '-0x2', '-0x1', '0x0', '0x3', '-0x1', '-0x2', '0x1', '0x0', '0x0', '0x1', '-0x1', '0x0', '0x2', '0x1', '-0x1', '-0x2', '-0x1', '-0x1', '0x1', '-0x1', '0x0', '0x0', '0x1', '0x1', '0x1', '0x0', '0x3', '0x0', '-0x1', '-0x3', '0x1', '-0x1', '0x1', '0x0', '0x2', '0x0', '0x2', '0x0', '0x1', '0x1', '0x1', '0x0', '-0x1', '0x0', '-0x1', '0x0', '-0x1', '0x1', '-0x3', '0x2', '0x1', '-0x1', '0x2', '-0x3', '0x2', '-0x2', '-0x1', '0x0', '-0x1', '0x1', '-0x1', '0x0', '0x1', '0x0', '0x0', '0x1', '-0x1', '0x1', '-0x1', '0x1', '0x1', '0x1', '0x1', '-0x1', '0x1', '-0x2', '0x0', '-0x2', '-0x1', '0x0', '0x1', '0x1', '-0x1', '-0x1', '-0x1', '0x1', '-0x1', '0x1', '0x0', '0x1', '0x1', '0x0', '0x2', '-0x1', '0x0', '-0x1', '0x1', '0x0', '0x1', '0x0', '0x2', '-0x1', '0x0', '0x0', '-0x2', '0x0', '0x1', '0x0', '-0x1', '-0x1', '0x0', '-0x2', '-0x1', '-0x1', '-0x2', '0x1', '-0x1', '0x0', '0x2', '0x1', '0x0', '0x2', '0x0', '-0x3', '0x0', '-0x1']
e
['-0x3', '0x2', '0x0', '0x0', '0x1', '0x0', '0x0', '0x0', '0x1', '-0x2', '0x0', '-0x1', '0x2', '0x1', '-0x2', '0x2', '0x0', '-0x2', '-0x1', '0x0', '0x0', '0x1', '0x1', '-0x1', '0x0', '0x0', '0x0', '0x1', '0x1', '0x1', '-0x1', '0x1', '0x1', '0x0', '-0x1', '0x0', '-0x1', '0x1', '-0x1', '-0x1', '0x0', '-0x1', '0x2', '0x3', '-0x2', '0x1', '0x1', '0x0', '0x2', '-0x1', '0x0', '-0x1', '0x1', '0x0', '-0x2', '0x2', '0x0', '-0x1', '0x0', '0x2', '0x0', '0x1', '-0x2', '0x0', '0x1', '0x1', '0x0', '-0x1', '-0x3', '0x0', '-0x1', '0x0', '-0x1', '0x1', '0x0', '0x1', '0x0', '0x1', '0x0', '0x1', '-0x1', '0x0', '-0x2', '0x2', '0x0', '-0x1', '-0x1', '0x0', '0x0', '0x1', '0x0', '0x1', '0x0', '-0x1', '-0x2', '0x0', '-0x1', '0x0', '0x0', '-0x1', '0x2', '0x0', '-0x1', '0x1', '-0x1', '-0x3', '-0x1', '-0x1', '0x1', '-0x1', '0x2', '0x1', '0x0', '0x0', '0x1', '0x0', '-0x1', '-0x1', '0x0', '0x0', '-0x1', '0x0', '0x3', '0x0', '0x1', '0x0', '0x1', '-0x2', '0x0', '-0x1', '0x1', '0x0', '0x0', '0x1', '-0x3', '0x0', '-0x2', '0x2', '0x0', '0x0', '0x0', '-0x1', '0x2', '0x0', '-0x1', '0x1', '0x2', '0x0', '0x0', '0x0', '-0x1', '0x2', '0x0', '0x0', '-0x1', '0x0', '-0x1', '0x0', '0x1', '0x0', '0x0', '0x0', '0x2', '-0x1', '-0x1', '-0x1', '-0x1', '0x2', '-0x1', '-0x1', '-0x1', '-0x1', '0x0', '-0x2', '0x1', '0x2', '-0x3', '0x2', '0x0', '0x2', '0x0', '0x0', '0x1', '0x1', '0x2', '0x0', '0x1', '-0x3', '0x1', '0x1', '0x2', '0x0', '0x3', '-0x2', '0x1', '0x2', '0x1', '0x0', '0x0', '-0x2', '-0x2', '-0x1', '0x0', '-0x1', '-0x3', '0x0', '0x1', '-0x1', '-0x2', '0x0', '0x1', '0x0', '0x1', '0x0', '-0x2', '-0x1', '0x0', '0x1', '-0x2', '0x0', '0x1', '0x1', '0x2', '-0x1', '-0x1', '0x2', '0x1', '-0x3', '0x2', '-0x2', '0x0', '-0x2', '0x0', '-0x1', '0x0', '0x1', '0x1', '0x1', '0x0', '0x0', '0x1', '0x1', '-0x1', '-0x1', '0x0', '-0x1', '-0x1', '-0x1', '-0x2', '0x0', '-0x1', '0x1', '0x0', '0x0', '0x0', '0x1']
['0x1', '0x0', '0x1', '-0x1', '0x0', '0x1', '0x0', '0x1', '0x2', '0x0', '0x0', '0x0', '0x1', '0x0', '-0x2', '0x1', '-0x1', '-0x1', '-0x1', '-0x2', '-0x2', '-0x1', '0x1', '0x0', '0x0', '0x0', '-0x2', '0x0', '0x0', '0x1', '0x1', '-0x3', '0x2', '0x0', '0x0', '0x0', '-0x1', '-0x2', '0x3', '-0x1', '0x0', '0x1', '0x0', '-0x1', '-0x1', '-0x2', '0x1', '0x1', '0x1', '-0x2', '0x0', '0x1', '-0x1', '-0x1', '-0x1', '0x1', '0x0', '0x1', '-0x1', '0x0', '0x1', '0x0', '0x1', '0x0', '-0x2', '0x0', '0x1', '0x1', '0x0', '-0x1', '0x0', '0x0', '0x1', '-0x1', '-0x2', '0x0', '-0x1', '0x1', '0x1', '0x1', '0x1', '-0x1', '0x2', '0x2', '0x0', '-0x1', '0x2', '0x2', '-0x2', '0x0', '0x1', '0x1', '0x3', '0x1', '0x0', '0x0', '-0x1', '0x2', '0x0', '0x2', '-0x2', '-0x1', '0x1', '-0x1', '0x0', '-0x1', '-0x1', '-0x1', '0x1', '0x0', '0x2', '-0x1', '0x1', '0x0', '0x1', '-0x1', '0x1', '0x0', '-0x1', '-0x1', '0x2', '0x2', '0x0', '0x3', '-0x2', '0x0', '0x2', '-0x1', '0x1', '0x0', '0x0', '0x0', '0x0', '0x0', '0x0', '0x0', '-0x2', '-0x3', '-0x3', '0x0', '0x0', '0x0', '-0x1', '0x1', '-0x2', '-0x1', '0x0', '0x1', '-0x2', '0x0', '-0x2', '-0x1', '0x1', '0x1', '0x2', '0x1', '0x1', '0x1', '0x0', '0x1', '0x0', '-0x2', '-0x1', '0x1', '-0x1', '-0x1', '0x0', '-0x1', '0x0', '0x0', '0x3', '-0x2', '0x0', '0x0', '0x0', '-0x1', '-0x1', '0x0', '0x3', '0x0', '0x1', '0x1', '-0x1', '-0x1', '0x0', '0x1', '0x0', '-0x1', '0x0', '0x1', '-0x1', '0x1', '0x2', '-0x1', '0x0', '0x1', '0x0', '0x1', '-0x1', '0x0', '-0x1', '0x0', '-0x1', '0x1', '-0x1', '0x1', '0x0', '0x3', '-0x1', '-0x1', '0x1', '0x0', '0x0', '0x0', '0x0', '0x2', '0x1', '-0x1', '0x1', '0x1', '-0x2', '0x1', '0x0', '0x0', '0x1', '0x3', '-0x1', '0x1', '0x3', '0x1', '0x0', '0x0', '0x1', '0x2', '0x0', '-0x2', '0x1', '0x0', '0x2', '0x0', '0x0', '0x0', '-0x2', '-0x1', '0x2', '0x1', '0x0', '-0x1', '0x0', '0x1', '0x0', '-0x2', '0x1', '0x1', '0x2', '-0x2']

*/