`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AIST
// Engineer: Junichi Sakamoto
// 
// Create Date: 2025/02/07
// Module Name: tb_sampler.sv
// Tool Versions: Vivado 2024.1
//////////////////////////////////////////////////////////////////////////////////



module tb_sampler;
    localparam integer
        CYCLE = 10,
        DELAY = 2,
        N_LOOP = 20;
                
    reg clk_i, rst_n_i, run_i;
    reg [255:0] rho_i;
    wire done_o;


    always begin
        #(CYCLE/2) clk_i <= ~clk_i;
    end

    sampleA dut(
        clk_i,
        rst_n_i,
        run_i,
        rho_i,
        done_o,
        polymat_A_o
    );

    /*-------------------------------------------
    Test
    -------------------------------------------*/
    initial begin
        clk_i <= 1;
        rst_n_i <= 1;
        #1000
        rst_n_i <= 0;
        run_i <= 0;
        rho_i <= reverse_endian_256(256'hc6195322bd2b71fd958cf071806587648fb31f7e4ee9ead48e0052b06244f3d1);
        #100
        rst_n_i <= 1;
        #5000;
        repeat (5) @(posedge clk_i);  // 5クロック後にrun_iを1にする
        run_i <= 1;
        repeat (1) @(posedge clk_i);  // 1クロック後にrun_iを0にする
        run_i <= 0;

        wait(done_o == 1);

        #1000
        rho_i <= reverse_endian_256(256'h7efb9e40c3bf0ff0432986ae4bc1a242ce9921aa9e22448819585dea308eb039);
        repeat (5) @(posedge clk_i);  // 5クロック後にrun_iを1にする
        run_i <= 1;
        repeat (1) @(posedge clk_i);  // 1クロック後にrun_iを0にする
        run_i <= 0;
    end

	function automatic logic [255:0] reverse_endian_256(input logic [255:0] data);
		logic [255:0] reversed = '0;

		for (int i = 0; i < 32; i++) begin
			reversed[i*8 +: 8] = data[(32-1-i)*8 +: 8];
    	end
    	return reversed;
	endfunction


endmodule

/*
For rho = 0xc6195322bd2b71fd958cf071806587648fb31f7e4ee9ead48e0052b06244f3d1

i=0,j=0
['0x456', '0x43c', '0x357', '0x9f4', '0x73f', '0x21c', '0xaa', '0x733', '0x135', '0xb5b', '0x43d', '0x543', '0x879', '0x5fe', '0x190', '0x715',
'0xc4c', '0x32', '0x701', '0x535', '0x9be', '0x622', '0x7be', '0xb24', '0x69f', '0x23', '0x59f', '0x961', '0xc89', '0xcbb', '0x278', '0x60',
'0x2a', '0xb68', '0x631', '0x738', '0x55f', '0x400', '0x314', '0x3b3', '0x860', '0x7ae', '0x61e', '0x712', '0x33b', '0x1e', '0x49e', '0x21e', 
'0xb18', '0x514', '0x7fc', '0x567', '0x850', '0x91d', '0xa27', '0x6a4', '0x4af', '0x6a9', '0xbc1', '0x1f0', '0xa0', '0x729', '0xb53', '0x73', 
'0x909', '0x7af', '0x8fa', '0xc99', '0x987', '0x47c', '0x567', '0x675', '0xc8c', '0x89', '0xb6', '0xa34', '0x8cc', '0xa36', '0x8fa', '0x453',
'0x62e', '0x4a5', '0x267', '0x531', '0x1d7', '0xc0b', '0xf5', '0x967', '0x96b', '0x2bc', '0xbf6', '0x14d', '0x9e7', '0x441', '0x520', '0x5aa',
'0xb91', '0x47a', '0x503', '0x7a4', '0x8f', '0x826', '0x695', '0x30a', '0x9f2', '0x903', '0xb6a', '0x72', '0x54', '0xcb2', '0xc4b', '0x39a', 
'0x7db', '0x8a0', '0x6b8', '0xb61', '0x5b4', '0xbe6', '0x549', '0x5be', '0x1b0', '0x568', '0x262', '0x8c1', '0x87', '0xa75', '0xa4b', '0x248', 
'0x23c', '0x126', '0x92', '0x764', '0x217', '0x959', '0x3b9', '0x277', '0x653', '0x770', '0xb08', '0x364', '0xadb', '0xa55', '0x528', '0x66d',
'0x946', '0x615', '0x304', '0x9d0', '0xb12', '0x492', '0x7d9', '0x9c6', '0x9c1', '0x76d', '0x282', '0x538', '0x32f', '0x75f', '0xb46', '0x1a3',
'0x7bc', '0x81a', '0x71a', '0x737', '0xbd3', '0x3c6', '0x6d1', '0x413', '0x76f', '0x61f', '0xb86', '0x6ad', '0xbfd', '0xccb', '0xc80', '0x338',
'0xbde', '0x97d', '0x7e0', '0x9a0', '0x348', '0x713', '0xa15', '0xac9', '0x9cc', '0x720', '0x801', '0xa3f', '0x90e', '0xb1d', '0x9d9', '0x5f3',
'0x1e9', '0x3fc', '0xabf', '0xab4', '0xcc3', '0x59b', '0x207', '0x12b', '0x970', '0x4c2', '0x9b4', '0xc53', '0x2dc', '0x9b5', '0xcf7', '0x2da', 
'0x324', '0xb9f', '0xa2e', '0x899', '0xbf3', '0x4f8', '0x3e9', '0xc75', '0x7e0', '0x5da', '0x529', '0xba0', '0x124', '0xadd', '0x276', '0xa90', 
'0x470', '0x97b', '0x68', '0x78c', '0x61e', '0x69d', '0x941', '0xafc', '0xac5', '0x150', '0x69c', '0xba4', '0x61b', '0x7cb', '0x1f5', '0x59a', 
'0x9fe', '0x651', '0x911', '0x6a7', '0x92d', '0x97b', '0x37a', '0x1e0', '0x743', '0x52f', '0x64', '0x2e7', '0x82f', '0xc01', '0xb50', '0x991']

i=0,j=1
['0x4ba', '0xb49', '0xab4', '0x729', '0x9c6', '0x291', '0xb48', '0xcc', '0xa1e', '0x820', '0x9ad', '0xdd', '0xb6c', '0x5fc', '0xbc9', '0x5', 
'0x397', '0x43e', '0xbdc', '0x866', '0x612', '0xa09', '0xcb6', '0xc77', '0xa27', '0x7f9', '0x408', '0xa60', '0x6e3', '0xc4a', '0x1a8', '0x9ec',
'0x631', '0x74e', '0x431', '0x6f4', '0x50d', '0xa03', '0x5d0', '0x8d3', '0x721', '0x620', '0x3e4', '0x322', '0x8da', '0x179', '0x206', '0xa97',
'0x436', '0x330', '0xa57', '0x4', '0x493', '0x470', '0xc5a', '0x361', '0x8c0', '0x831', '0xabb', '0xf4', '0x78', '0x3f9', '0x58e', '0x2d6',
'0x21c', '0x66e', '0x3d6', '0x21a', '0x37b', '0xc7a', '0x5f4', '0x168', '0xb12', '0x91', '0x1d7', '0x529', '0x363', '0xba1', '0x5c2', '0x10e',
'0x1dc', '0x5f3', '0x110', '0xbe1', '0x16b', '0xcd1', '0x5af', '0x891', '0x26b', '0x35', '0xb62', '0x861', '0xa25', '0x980', '0x3e7', '0x571', 
'0xfb', '0x8fb', '0x92d', '0x717', '0x3e6', '0x717', '0x877', '0x2b2', '0x819', '0x988', '0x527', '0xba9', '0x4e9', '0x19', '0x46c', '0x422',
'0x392', '0x503', '0x974', '0x2c3', '0x757', '0x3d4', '0xa9', '0x45b', '0x79c', '0x916', '0x25', '0xa2f', '0x7e8', '0x4b5', '0x2cf', '0x840',
'0x3d9', '0xa88', '0x7d7', '0xb22', '0x591', '0x67a', '0xc1c', '0xc3', '0x92b', '0x3af', '0xbcf', '0xa38', '0x74c', '0x8bd', '0xbc', '0x9be',
'0x99', '0x7dc', '0x5d', '0xb69', '0xcc8', '0x80f', '0xb71', '0x9ef', '0x9c4', '0xae4', '0x3d7', '0x5b7', '0x557', '0x3f6', '0x137', '0x7e6',
'0xb92', '0x641', '0x3a6', '0x3a2', '0xa1a', '0x5cd', '0x34f', '0xa02', '0x27f', '0xb9f', '0x7f7', '0x952', '0xc59', '0x800', '0x604', '0xc',
'0x19f', '0x57f', '0x46', '0x6f0', '0x655', '0xc3f', '0x4b1', '0x726', '0x242', '0x814', '0xa88', '0x59b', '0xa3b', '0xb41', '0xb3f', '0xc92',
'0x213', '0x5e0', '0x8ca', '0x69a', '0x2b5', '0x972', '0x742', '0xa72', '0xb35', '0xb76', '0xcb8', '0x881', '0x4b3', '0x2b2', '0x416', '0x396', 
'0x34f', '0x9c5', '0x521', '0xcfe', '0x5ec', '0x310', '0x48d', '0x6e3', '0x72b', '0xbd7', '0x748', '0x811', '0xb3b', '0x6a9', '0xabd', '0x825',
'0x487', '0x38d', '0xb8', '0xc92', '0x6e0', '0x709', '0x95', '0x2c', '0x1e6', '0x82b', '0x6fc', '0x29', '0x842', '0x1cc', '0x739', '0x713',
'0x703', '0xcf3', '0x1ae', '0x70e', '0x7c', '0xcf2', '0x294', '0x393', '0x489', '0xa61', '0x29a', '0x940', '0xcb4', '0x10', '0x908', '0x77']

i=1,j=0
['0x690', '0x416', '0x136', '0x882', '0x77a', '0x937', '0x61f', '0xcc9', '0xcdc', '0x5f4', '0x927', '0xaa0', '0x2e', '0x602', '0x992', '0xe8', '0x625', '0xadd', '0x276', '0x645', '0x6c5', '0x5b6', '0x9a', '0xc05', '0xc73', '0x393', '0x631', '0x365', '0x794', '0x319', '0x27b', '0x4ef', '0xa99', '0x435', '0x172', '0x5c2', '0x32f', '0x8c6', '0x934', '0x8ae', '0x2b5', '0x4e2', '0xbbd', '0x5c8', '0xbca', '0x2cd', '0x35c', '0xcf7', '0x80c', '0xb88', '0xa18', '0x9ad', '0xbcf', '0x88b', '0x558', '0x59', '0x800', '0x51e', '0x6b2', '0x11e', '0x660', '0x4b1', '0x6ea', '0x81a', '0x1e', '0xbf6', '0xa83', '0xc42', '0x94f', '0xa2c', '0x730', '0x2fd', '0xa00', '0xb08', '0xbd9', '0x1de', '0x93a', '0x43c', '0x3fd', '0x7ba', '0xca9', '0xccc', '0x83', '0x87c', '0xc90', '0xb25', '0x5de', '0x831', '0x54c', '0x95d', '0x560', '0xbc', '0x55', '0x841', '0x61f', '0x848', '0x959', '0x30c', '0x98e', '0x716', '0xc1d', '0x3e8', '0x726', '0x524', '0x923', '0x7e0', '0x3e7', '0x709', '0x1d3', '0x21a', '0xc68', '0xabb', '0x82b', '0xc01', '0x4c3', '0x4e8', '0xf4', '0xc71', '0x597', '0xce9', '0x3c4', '0xc84', '0x638', '0xa68', '0xc6', '0x3a3', '0xc1c', '0x967', '0xabc', '0x703', '0xa60', '0x7a1', '0x210', '0x857', '0x933', '0x697', '0x32c', '0x17b', '0x1c6', '0x6ab', '0x6ab', '0x501', '0xabb', '0x512', '0x31', '0xe3', '0x578', '0xbbd', '0x3d8', '0xb93', '0xaa4', '0x199', '0xbc2', '0x24b', '0x93c', '0x840', '0x6b5', '0x627', '0xaa0', '0x318', '0x8c', '0x8d6', '0x5d1', '0x3bb', '0xf7', '0x7da', '0x453', '0x824', '0x855', '0x1a', '0x6d8', '0x37d', '0x84a', '0x3d', '0x654', '0x251', '0x78a', '0xc8', '0x1ba', '0x6dc', '0x91a', '0x326', '0x654', '0x6c4', '0xac', '0x83c', '0x33', '0xa23', '0x6e9', '0x5c1', '0x74f', '0x5b7', '0x3fd', '0x8c0', '0xa7a', '0xcb7', '0xabc', '0x552', '0x6fb', '0x697', '0x6a2', '0x890', '0x601', '0xcb0', '0x1ad', '0xbe', '0x83', '0x6fd', '0x977', '0x58c', '0x538', '0x72e', '0x5c4', '0x72b', '0x573', '0x5d2', '0x2a2', '0x231', '0xae0', '0x3d2', '0x3ed', '0xb8d', '0xae7', '0x4ce', '0x7ca', '0x4d7', '0x17c', '0x282', '0x626', '0x30', '0x112', '0xa8b', '0x79c', '0x634', '0x39a', '0x87c', '0xc6b', '0x562', '0x5d2', '0x406', '0xbd4', '0xa9b', '0xcf5', '0x4fc', '0x214', '0x89b', '0x97f', '0xc49', '0x748', '0x66a', '0xbce', '0xa', '0x8fc', '0x7b8', '0x82', '0x9b2']

i=1,j=1
['0x5e1', '0x336', '0xc7f', '0xabf', '0x4fc', '0x682', '0x495', '0x9fd', '0x23d', '0x69', '0x1e1', '0x5d3', '0x539', '0x698', '0x3f0', '0x305', '0x6e7', '0xa8e', '0x5e0', '0x630', '0xb8b', '0x4e9', '0x9ad', '0x8fb', '0x1dc', '0x400', '0x37d', '0xc5d', '0x199', '0xf8', '0x505', '0x5e3', '0x5e0', '0x7e', '0x690', '0x6b3', '0x9b6', '0x977', '0x1e', '0x209', '0xbdd', '0x48a', '0x64f', '0xa19', '0x591', '0x2ad', '0xc9a', '0x415', '0x29a', '0x967', '0xa34', '0x345', '0x69d', '0x1bb', '0x66c', '0x5d3', '0x8b9', '0x332', '0x576', '0x3f8', '0x645', '0x7be', '0xbc4', '0x93f', '0x5f9', '0x450', '0x130', '0x17c', '0xbde', '0x9af', '0xa7e', '0x969', '0x7e3', '0xc4d', '0x9f8', '0x5ef', '0x35', '0xcf7', '0x51f', '0xa51', '0x7b3', '0x243', '0x4f5', '0x34b', '0x23e', '0x480', '0x924', '0xcb7', '0x5b3', '0xa', '0x69b', '0x188', '0x117', '0x9e8', '0x8bc', '0xa99', '0x7d1', '0x2f9', '0xc10', '0x2c0', '0x11b', '0x7b0', '0x857', '0x792', '0x32b', '0x26f', '0x7f7', '0x5df', '0xf3', '0x591', '0x394', '0x39c', '0xacf', '0xb2a', '0x57e', '0xf9', '0x239', '0x76', '0x6af', '0xbe9', '0x1ae', '0x78b', '0x126', '0x358', '0x350', '0x25a', '0x924', '0x48f', '0xbaf', '0x10d', '0x378', '0x941', '0x11', '0x1b5', '0x532', '0x7ac', '0x599', '0x384', '0xaf', '0x9c6', '0xc88', '0xc6a', '0x1e', '0xb78', '0x990', '0x6c3', '0x90', '0xb31', '0x38b', '0x1fa', '0x9e8', '0x9b4', '0x1f2', '0xb63', '0xbfd', '0x19c', '0xb49', '0x10a', '0x671', '0x624', '0xc62', '0xb43', '0x19a', '0x14d', '0xb75', '0x8d6', '0xca5', '0x363', '0x7cc', '0x5b8', '0x340', '0xc27', '0x303', '0xc0a', '0x26d', '0x639', '0x3a', '0x9db', '0x932', '0x610', '0x8cb', '0xb6e', '0xc54', '0x182', '0x29d', '0xaee', '0x431', '0x15', '0x985', '0x616', '0x9ef', '0x87a', '0x872', '0x938', '0x76', '0x50d', '0x29c', '0x9', '0xb9f', '0x2a7', '0x88', '0x41', '0xad7', '0xc8a', '0x1dc', '0x4ef', '0x89b', '0xce5', '0x96e', '0x738', '0xb9a', '0x58d', '0x225', '0xc59', '0x2bb', '0x289', '0xa78', '0x895', '0xc80', '0x2bc', '0xb6a', '0xaa9', '0x56', '0x782', '0x2ed', '0xadf', '0x2', '0x5b5', '0xcf5', '0x2c7', '0x576', '0x2a5', '0x5f3', '0xbed', '0x5b5', '0x52e', '0x79', '0xa12', '0x5c9', '0x1a', '0x957', '0x4c4', '0x29f', '0x919', '0x824', '0x912', '0x124', '0x30c', '0x328', '0x581', '0x5aa', '0x97a', '0xac1', '0xcda', '0x6a6', '0x675']


For rho = 0x7efb9e40c3bf0ff0432986ae4bc1a242ce9921aa9e22448819585dea308eb039

['0x5a9', '0xabc', '0x50f', '0x45f', '0x168', '0xbca', '0xa4b', '0xb7e', '0x663', '0x77e', '0x12f', '0x7b4', '0x409', '0x164', '0x75f', '0x409', '0xc65', '0x307', '0x567', '0x609', '0x707', '0xa1c', '0x17', '0x8fe', '0x99d', '0xac3', '0x75', '0x95a', '0x106', '0x22f', '0x406', '0x946', '0x7b7', '0x847', '0x815', '0x667', '0x407', '0x466', '0x352', '0x83e', '0x833', '0x478', '0xc3d', '0x6d7', '0x61d', '0x3fa', '0x85', '0x682', '0x417', '0x278', '0xc29', '0x54b', '0x757', '0xcb0', '0x2de', '0x469', '0x1a6', '0x972', '0xb06', '0x77d', '0xcf4', '0x8c', '0x5c', '0x1eb', '0x97a', '0x164', '0x81f', '0x9a1', '0x804', '0xa2e', '0xc21', '0x379', '0x7be', '0x830', '0xb58', '0x2fb', '0xe7', '0x994', '0xaa1', '0x487', '0xcfb', '0x6eb', '0x844', '0x90d', '0xa71', '0x418', '0xbb5', '0xadd', '0x938', '0x2da', '0xbd9', '0x52a', '0x7a6', '0x74f', '0x240', '0xbab', '0x6fd', '0x735', '0xd00', '0x699', '0x8b7', '0x194', '0xc11', '0xc1', '0x807', '0x60b', '0x3cf', '0x461', '0x467', '0x46d', '0x480', '0xcea', '0xa48', '0xa4f', '0x57e', '0xc7d', '0x9de', '0x82', '0xb31', '0x1d2', '0x1b4', '0x9a9', '0x4bb', '0xc19', '0xc7f', '0xcf9', '0xc03', '0x9cb', '0x4ad', '0x68c', '0xf7', '0x9ab', '0x25c', '0xadb', '0x88', '0xad0', '0x192', '0x273', '0x53d', '0xa24', '0x1ea', '0x346', '0xc79', '0x27', '0x84b', '0x80f', '0x329', '0x2e1', '0x816', '0x26e', '0x610', '0x17f', '0x916', '0x3b8', '0x61b', '0x20e', '0x6bd', '0xb76', '0x57b', '0x336', '0x42c', '0x3ad', '0xc25', '0x66e', '0x1b4', '0x942', '0x615', '0xca2', '0x4c0', '0x9a6', '0x23c', '0x509', '0xf7', '0x95a', '0x17c', '0x3b1', '0x5dc', '0x84d', '0xa92', '0x668', '0x976', '0xb71', '0x17e', '0x30d', '0x81b', '0xb19', '0x3d6', '0xa21', '0x30', '0x9ec', '0x1ad', '0xae3', '0x66f', '0x27f', '0x7a5', '0x270', '0x489', '0x38c', '0xa93', '0x4be', '0x8fc', '0x99', '0x81a', '0xc33', '0xa2', '0x19b', '0xb76', '0xc5c', '0x44', '0x3d6', '0x69d', '0x810', '0x70e', '0x1b0', '0xc8f', '0xc8b', '0x44c', '0xa32', '0x58', '0xc9d', '0x1a5', '0x6b7', '0x3ac', '0x12e', '0x4a9', '0xcf', '0xc8a', '0x2d4', '0xb06', '0xb07', '0x856', '0x8b6', '0x52e', '0xb3f', '0xb40', '0x651', '0x727', '0xae9', '0x92b', '0x17', '0xa66', '0x11e', '0x245', '0x115', '0x42d', '0x7c', '0xd2', '0xc72', '0xb67', '0xba1', '0x931', '0x810', '0x1ad', '0x7bc', '0x449', '0xc0']

['0xa3b', '0x223', '0x9ba', '0x841', '0xd3', '0x5b2', '0x8ce', '0x408', '0x12c', '0x986', '0xaf3', '0x652', '0x895', '0xcef', '0x7b3', '0x445', '0x592', '0x829', '0x6b0', '0x421', '0x81f', '0x4d6', '0x23f', '0x842', '0x79b', '0xafb', '0x5c9', '0x3dc', '0x4c9', '0x63a', '0x587', '0x7ad', '0x3f', '0x8', '0x1f', '0x19', '0xc92', '0xcd6', '0xa44', '0x2c', '0x56f', '0x8dc', '0x25f', '0x8cf', '0x97f', '0x3b3', '0xa0a', '0x473', '0x19e', '0x8df', '0x775', '0x8f1', '0x4f', '0xc4b', '0x8e1', '0x736', '0x846', '0x3a8', '0xc48', '0x4e8', '0x2a9', '0x518', '0xa6f', '0x51a', '0xa66', '0x597', '0xb8', '0xce8', '0x360', '0xbf6', '0x607', '0x241', '0x130', '0x81a', '0x1ce', '0xb77', '0x420', '0xc9e', '0x28a', '0x3f1', '0x58d', '0x7ca', '0x766', '0x646', '0x423', '0x51b', '0x4b8', '0x184', '0xdb', '0xd2', '0x152', '0x87d', '0x346', '0x4f7', '0xcf6', '0x44e', '0x7d4', '0xb79', '0xa32', '0x766', '0x60d', '0xc27', '0x5db', '0xa06', '0x876', '0x79a', '0x266', '0xf3', '0x42', '0x8f', '0x2a9', '0x63e', '0x720', '0xabf', '0xc01', '0x3dc', '0x9b5', '0xe0', '0x41b', '0x462', '0x110', '0xd2', '0xa22', '0x7ec', '0xa1d', '0x13f', '0x852', '0x947', '0xbee', '0xbbf', '0x1ef', '0x933', '0x1e5', '0x3cb', '0x7a9', '0x9af', '0xaaf', '0xa5c', '0x25', '0x661', '0x449', '0x52a', '0xc7', '0xa6e', '0x7fd', '0xb53', '0x779', '0x6cc', '0xa35', '0x3a', '0xbe7', '0x919', '0x89', '0xbf0', '0x5e1', '0xa86', '0x1d', '0x17d', '0xaaf', '0x649', '0x4a0', '0x16c', '0x505', '0x75e', '0x67a', '0xcda', '0x48e', '0x6d', '0x787', '0x92e', '0x380', '0x1cf', '0x93c', '0x1cb', '0x1c0', '0xbcc', '0x2b4', '0x590', '0x680', '0x3b', '0x56a', '0x534', '0xb49', '0x41e', '0x4a8', '0x76e', '0x9b8', '0x93e', '0x281', '0x263', '0xa50', '0x4e4', '0xaeb', '0x8ac', '0xbde', '0xc27', '0xabb', '0x8a5', '0xbf9', '0x8db', '0xaec', '0x212', '0x65c', '0x986', '0x3a8', '0xc60', '0x197', '0xbb', '0x870', '0xe9', '0x7dc', '0x925', '0x3bd', '0x344', '0x46d', '0x1b3', '0x1d8', '0x7bd', '0x702', '0x585', '0x5c9', '0xaa4', '0x5', '0xaaf', '0x35d', '0x6c8', '0xbd2', '0x86a', '0x6c6', '0x14b', '0xb3d', '0x58', '0xb7b', '0x916', '0x4c6', '0x9d5', '0xad5', '0xb0f', '0x41c', '0x868', '0x78c', '0x3ce', '0x568', '0x10', '0x7a6', '0xc01', '0x606', '0x70a', '0x1e6', '0x583', '0xc7f', '0x571', '0x244', '0xc4d', '0x8b1', '0x6dd']

['0x22e', '0x81e', '0x5f9', '0x128', '0x7cc', '0x5c1', '0x60a', '0x1d', '0x6d', '0x83', '0x478', '0x9e6', '0x21c', '0xcbe', '0x442', '0xc48', '0xb48', '0xa3e', '0x7df', '0x3a4', '0x911', '0x3a5', '0x47a', '0x517', '0x43a', '0xc6e', '0xbab', '0x19b', '0xca5', '0x649', '0xae8', '0x718', '0xce4', '0xbaf', '0x14', '0x5a8', '0x1b4', '0xb83', '0x7c7', '0x24b', '0xb9c', '0xba9', '0x65', '0xc1a', '0x4cb', '0x4b9', '0x8f5', '0xa0a', '0x623', '0x12a', '0x7f1', '0x733', '0xbd', '0x472', '0xc57', '0x941', '0x7b4', '0x66e', '0x3e6', '0x895', '0x83', '0x432', '0x3df', '0x9a1', '0x68c', '0x964', '0xa58', '0x947', '0xbd9', '0xc66', '0x238', '0x2fc', '0x5cc', '0x1f1', '0xa43', '0x8f1', '0x3af', '0xa62', '0x922', '0xa8f', '0x4cc', '0xb00', '0x12b', '0x12b', '0x5ad', '0xad9', '0x628', '0xb3d', '0x2c1', '0xb85', '0x930', '0x57e', '0xc3f', '0x668', '0x2a1', '0xcfb', '0xcfa', '0x1fe', '0x3b4', '0xf7', '0xbb1', '0xc10', '0x562', '0x86d', '0x152', '0xc6d', '0xca4', '0x280', '0xc44', '0xa94', '0x8e4', '0xab5', '0x294', '0xa4d', '0xb7a', '0x294', '0xb4e', '0xa45', '0x2a5', '0x2c9', '0x16b', '0xa98', '0x709', '0x12b', '0x19c', '0xc7d', '0x571', '0x81d', '0xa97', '0x5a5', '0x71', '0x4fa', '0x8d8', '0x2f3', '0x7f6', '0x650', '0x423', '0x710', '0xbf6', '0xb27', '0x546', '0x89', '0xcaf', '0xb7', '0x520', '0xa3a', '0x13', '0x54d', '0xb14', '0x842', '0x7c4', '0xc7', '0x370', '0x958', '0x6ff', '0x1b2', '0x457', '0x58', '0x7b1', '0x71f', '0x9a4', '0x372', '0x59f', '0xb5f', '0xc7b', '0x1c1', '0xe4', '0x15f', '0x355', '0xb5c', '0x89f', '0x839', '0x86a', '0xbe0', '0x5fc', '0x69d', '0x1ec', '0x286', '0x130', '0x527', '0xafe', '0x4c7', '0x79e', '0xd7', '0x97', '0x992', '0x75a', '0xaae', '0x555', '0x98e', '0xc21', '0xb93', '0xb8d', '0x9b6', '0x400', '0xa66', '0x2fd', '0xc6b', '0x81b', '0x981', '0x763', '0x2c1', '0xbf2', '0xc5a', '0xce9', '0x37c', '0x72e', '0x3a3', '0x670', '0x593', '0x264', '0x410', '0x2d9', '0x9e8', '0x2f', '0x20f', '0xbdf', '0xbb5', '0x9ab', '0xadd', '0x7d7', '0xca4', '0x7ed', '0xbd0', '0x339', '0x8dc', '0x185', '0x151', '0x327', '0x691', '0x410', '0x43c', '0x99c', '0x6a9', '0xaaf', '0x38', '0x2dd', '0x844', '0x82f', '0xa0f', '0x14', '0xcbb', '0x26e', '0x5a7', '0xc55', '0xb09', '0xc22', '0xae2', '0xb80', '0x912', '0x454', '0xc84', '0x2c2', '0x7d4', '0xc9d', '0xb98']

['0x653', '0x4e', '0x775', '0x5b6', '0xb34', '0xbb8', '0x475', '0x2cd', '0x103', '0x72c', '0xbdd', '0xcac', '0xca', '0xca0', '0x7f2', '0x214', '0xbfe', '0x771', '0x74d', '0x45a', '0xaae', '0x487', '0x146', '0x902', '0x5a0', '0xb36', '0x690', '0xb47', '0x29a', '0x12e', '0x3e4', '0x92e', '0x585', '0x79b', '0x684', '0x371', '0x80c', '0xc64', '0x49f', '0xa2c', '0x4', '0x36f', '0xaec', '0x418', '0xbe1', '0x2bd', '0xd00', '0x827', '0x216', '0x988', '0x33a', '0x4d5', '0xc08', '0x49e', '0xc7', '0x65d', '0x84a', '0x8e4', '0xb87', '0x9eb', '0xe5', '0x1f8', '0x9c1', '0x3f3', '0x4da', '0x239', '0xacb', '0x8af', '0x40b', '0x903', '0x8ab', '0x510', '0x305', '0xc82', '0xa18', '0x4c1', '0x8a6', '0x34f', '0xb5f', '0xa89', '0x88f', '0xc0c', '0xc65', '0xb53', '0x361', '0x9a', '0xa67', '0x8d2', '0x7fa', '0x676', '0x750', '0xcbf', '0x9c3', '0x57c', '0xa5c', '0x283', '0x5da', '0xb63', '0x824', '0xbc5', '0x4a4', '0x4ba', '0xa6f', '0x28b', '0xb78', '0x8bd', '0x810', '0x80c', '0x46e', '0xbc6', '0xc9e', '0xf6', '0x893', '0xab0', '0x99c', '0xcd', '0xc2a', '0x231', '0x78a', '0x648', '0xa9', '0x98f', '0x3e0', '0x733', '0x5ea', '0xfc', '0x8ee', '0x29', '0x3c6', '0x136', '0x209', '0x170', '0xac4', '0x912', '0xb41', '0xbb5', '0x32a', '0x1db', '0x6a7', '0x4e', '0x45d', '0x2f2', '0xcff', '0x277', '0x534', '0x2f8', '0x35a', '0x99e', '0xe5', '0x913', '0xcfe', '0x916', '0x5cf', '0x8cf', '0x22c', '0x5fa', '0x2fe', '0x88f', '0xc95', '0x934', '0x3f7', '0xad2', '0xb69', '0x489', '0x9cb', '0x34e', '0x15a', '0x800', '0x800', '0x888', '0x2be', '0x947', '0x9e8', '0x776', '0x7a3', '0x1fa', '0x9af', '0x935', '0x889', '0x220', '0x9d7', '0xcc1', '0x997', '0x17d', '0x231', '0xb', '0x60a', '0x408', '0x103', '0x62c', '0x962', '0x62a', '0x612', '0x392', '0x572', '0x4f1', '0x792', '0x1da', '0x8f4', '0x26d', '0xc5c', '0x185', '0x39', '0x3b9', '0x1cb', '0xb8c', '0xc06', '0xba3', '0x52', '0x5d0', '0x104', '0x70a', '0x161', '0x2d7', '0xb2d', '0x277', '0x4da', '0x66e', '0x797', '0x148', '0x72e', '0xa75', '0xc98', '0x406', '0x838', '0x192', '0x8fd', '0xbe5', '0x556', '0x357', '0x54b', '0x9f9', '0x2aa', '0x713', '0xb06', '0x8be', '0xaaa', '0x1e', '0xb2', '0x3ed', '0x6dc', '0x8c1', '0x511', '0x692', '0x1bb', '0xc98', '0x411', '0xbc4', '0x7e7', '0xca7', '0x8ae', '0xcf2', '0x77f', '0xc1e', '0xb5e', '0x2c5']

*/

