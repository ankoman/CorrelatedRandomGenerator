`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AIST
// Engineer: Junichi Sakamoto
// 
// Create Date: 2024/02/05
// Module Name: sampleA
// Target Devices: U250
// Tool Versions: Vivado 2024.1
//////////////////////////////////////////////////////////////////////////////////


module sampleA
     import TYPES_KEM::*;
    (
        input clk_i,
        input rst_n_i,
        input run_i,
        input [255:0] rho_i,
        output done_o,
        output polymat_t polymat_A_o
    );
    localparam CNT_WIDTH = $clog2(ML_KEM_K*ML_KEM_K);
    localparam K_WIDTH = $clog2(ML_KEM_K);


    logic [CNT_WIDTH:0] cnt_kk;
    wire sample_run, sample_rdy, sample_done, busy;
    logic [K_WIDTH - 1:0] index_i, index_j;
    poly_t poly_o;

    assign busy = |cnt_kk;
    assign sample_run = run_i || (sample_done && busy);
    assign sample_done = done_o;
    assign done_o = cnt_kk[CNT_WIDTH] && sample_done; // ML-KEM-512 specific definition
    assign index_i = cnt_kk[0]; // ML-KEM-512 specific definition
    assign index_j = cnt_kk[1]; // ML-KEM-512 specific definition

    always_ff @(posedge clk_i) begin
        if(!rst_n_i || done_o) begin
            cnt_kk <= '0;
        end
        else if(sample_run) begin
            cnt_kk <= cnt_kk + 1'b1;
        end
    end

    sampleNTT u0(
        .clk_i,
        .rst_n_i,
        .run_i(sample_run),
        .rho_i,
        .index_i_i(8'(index_i)),
        .index_j_i(8'(index_j)),
        .done_o(sample_rdy),
        .poly_o
    );

    always_ff @(posedge clk_i) begin
        if(!rst_n_i)
            polymat_A_o <= '0;
        else if (sample_done)
            polymat_A_o[index_j][index_i] <= poly_o;
    end

endmodule

module sampleNTT
     import TYPES_KEM::*;
    (
        input clk_i,
        input rst_n_i,
        input run_i,
        input [255:0] rho_i,
        input [7:0] index_i_i,
        input [7:0] index_j_i,
        output done_o,
        output poly_t poly_o
    );

    keccak_1600_t xof_in, xof_out;
    logic [4:0][63:0] xof_msg;
    assign xof_msg = {40'd0, 8'h1f, index_i_i, index_j_i, rho_i};

    assign xof_in[0][0] = xof_msg[0]; // [63:0]
    assign xof_in[1][0] = xof_msg[1]; // [127:64]
    assign xof_in[2][0] = xof_msg[2]; // [191:128]
    assign xof_in[3][0] = xof_msg[3]; // [255:192]
    assign xof_in[4][0] = xof_msg[4]; // [319:256]
	assign xof_in[0][4] = 64'h8000000000000000;
    generate
        for(genvar i = 1; i < 5; i = i + 1) begin
            for (genvar j = 0; j < 5; j = j + 1) begin
                if((i == 4) && (j == 0)) begin
                    // Do nothing
                end
                else
                    assign xof_in[j][i] = 64'h0;
            end
        end
    endgenerate

    logic xof_rdy, xof_rdy_prev;
    logic [6:0] cnt_112;
    logic [7:0] cnt_sampled_coeff, cnt_squeezed;
    logic [1343:0] xof_rate;
    wire xof_run = run_i | sample_end;

    always_ff @(posedge clk_i) begin
        xof_rdy_prev <= xof_rdy;
    end
    wire sample_start = ({xof_rdy_prev, xof_rdy} == 2'b01) ? 1'b1 : 1'b0; // Rising edge. Same time as squeeze done.
    wire sample_end = (cnt_112 == 7'd112) ? 1'b1 : 1'b0;
    wire sample_busy = |cnt_112;
    wire [ML_KEM_LEN_Q - 1:0] coeff = xof_rate[ML_KEM_LEN_Q - 1:0];
    wire is_reject = (coeff > (ML_KEM_Q - 1)) ? 1'b1 : 1'b0;
    wire sel_xor_in = |cnt_squeezed;
    assign done_o = (cnt_sampled_coeff == 8'hff);

    always_ff @(posedge clk_i) begin
        if(!rst_n_i | done_o) begin
            cnt_squeezed <= '0;
        end
        else if(xof_run) begin
            cnt_squeezed <= cnt_squeezed + 1'b1;    // If overflowing, then should abort
        end
    end

    always_ff @(posedge clk_i) begin
        if(!rst_n_i || sample_end || done_o) begin
            cnt_112 <= '0;
        end
        else if(sample_start | sample_busy) begin
            cnt_112 <= cnt_112 + 1'b1;
        end
    end

    always_ff @(posedge clk_i) begin
        if(!rst_n_i || done_o) begin
            poly_o <= '0;
            cnt_sampled_coeff <= '0;
        end
        else if(sample_busy && !is_reject) begin
            poly_o <= {coeff, poly_o[255:1]};
            cnt_sampled_coeff <= cnt_sampled_coeff + 1'b1;
        end
    end

    always_ff @(posedge clk_i) begin
        if(!rst_n_i) begin
            xof_rate <= '0;
        end
        else if(sample_start) begin
            xof_rate <= xof_out[1343:0];
        end
        else if(sample_busy) begin
            xof_rate <= {12'd0, xof_rate[1343:12]};
        end
    end

	keccak_top #(.d(0), .b(1600), .W(64)) xof (
		.Clock(clk_i), 
		.Reset((!rst_n_i) | xof_run), 
		.InData(sel_xor_in ? xof_out : xof_in), 
		.FreshRand(), 
		.Ready(xof_rdy), 
		.OutData(xof_out)
	);

endmodule
