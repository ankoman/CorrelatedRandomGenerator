`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AIST
// Engineer: Junichi Sakamoto
// 
// Create Date: 2024/10/26
// Module Name: test_aes.sv
// Tool Versions: Vivado 2020.1
//////////////////////////////////////////////////////////////////////////////////



module test_aes_uart;
    localparam 
        CYCLE = 10,
        DELAY = 2,
        N_LOOP = 20;
                
    reg clk, rst_n, uart_rx;
    reg [23:0] cycle_cnt;

    always begin
        #(CYCLE/2) clk <= ~clk;
    end

    TOP_CRG_HW_UART dut(
        .CLK100MHZ(clk),
        .ck_rst_n(rst_n),
        .uart_txd_in(uart_rx),
        .uart_rxd_out(),
        .led()
    );

    /*-------------------------------------------
    Test
    -------------------------------------------*/
    initial begin
        clk <= 1;
        rst_n <= 1;
        #1000
        rst_n <= 0;
        uart_rx <= 1;
        #100
        rst_n <= 1;
        #1000;
        UART_RX_128(8'h10, 8'h00, 128'h2b7e151628aed2a6abf7158809cf4f3c);   // Set key
        #1000
        UART_RX(8'h40);  // Run
        #1000
        $finish;
    end

    task UART_RX;
        parameter   RATE=115200;//ボーレート[bps]
        input[7:0]  dat;//送るデータ  
        integer     i;//ループ用変数
        time        BIT_CYC;//1ビットの周期
    
        begin
            $display("UART input start : 0x%2X",dat);
            //ボーレートからbit周期[ns]を算出
            BIT_CYC=1000000000/RATE;//timescaleが1nsの前提
            //スタートビット
            uart_rx  <=1'b0;
            #BIT_CYC;
            //データ:LSBファースト
            for(i=0; i<8; i=i+1)begin
                uart_rx <= dat[i];
                #BIT_CYC;
            end
            //ストップビット
            uart_rx <= 1'b1;
            #BIT_CYC;
        end
    endtask

    task UART_RX_128;
        integer i;
        input [7:0] com;
        input [7:0] addr;
        input [127:0] dat;
        
        begin
            UART_RX(com);
            UART_RX(addr);
            for(i = 0; i < 16; i=i+1) begin
                UART_RX(dat[7:0]);
                dat = {8'd0, dat[127:8]};
                #1000;
            end
        end
    endtask

endmodule

/////////////////////////////////////////////////////////////////////
// PRNG256 Test vectors, key = 0x2b7e151628aed2a6abf7158809cf4f3c
/////////////////////////////////////////////////////////////////////
// 0x7df76b0c1ab899b33e42f047b91b546ff6c71eedc3d99bb183cb5b8d1568e606
// 0x57127d4034b1bebfaef466b9c7726fc633d495111a4b3d37cc76f29c3398894f
// 0x973f2ef34879e2027f1734303ff21f894106dc419a06db149dd22bfb583ffeee
// 0x469c7fcb75d5d9a1b418cb997b09a185e2c75fad134f621d9223df0a9c2793d8
// 0x8a7c37ad7c3edf32495ececadec2311cd39847fd634a2b73f776242e3dedcf1f
// 0xef28d82739fd8c7147323f7e91c0cbface3030cf459b183beaf59fed49fa8d10
// 0x3066e41e679d88b8efeb7b3d4af3f6c1345fc1e3ba0123d0024cd00b579e7b01
// 0x8b6af01acb7464cb68c4a3548aaf95a67784d2a5aac5066e710a151d5590c008
// 0xc7ca47a1df471b5a273fec3be2e595bb936ce9493f3a5c5d720798aaa3f77a3
// 0x3f73d097873e5a3ef789572193bb63a250563c6b25399ca756e342bd24eb2ec3
// 0x71577831908d0b644c364131acfb0a63613f5a9ff21cb9f251990f54e5669168
// 0xd3ccd84141e0772ac5ff9995184621f4d714c1895acf07d243f64cd232780bd5
// 0xf201fa2e105087f23751f7f586b430d36bd47571e4d5ab2570ee08cdd1c36773
// 0x1f39117775381545539d17d6872a28b1d60250445609c944dcd632c561d12cea
// 0x861c5964e3c9dc95c6303f12bad10d9c424cb3cbe88e15c8844be3802d5f3dcc
// 0x53274720b085c306d508e9fd7928624fef6be65d9a0da57aefd277cfb4a06e66
// 0x7e794a13c74973b4bf55b10f5a9904e85d292b7950100926cab2d1313937b41d
// 0x46440182b842e3af60292498ea18ea42bc94af882df59e87a8572648cd769a4c
// 0x20c4647cd97571b5b142b8ea289619e0a8b50c49f12b034827d3e5c1580352ef
// 0x3afb2a4eb995fda13ff080b05eae6cfdf3464517146d3a60946197e455fe69a3
// 0x56980cee98e1b9b47a0f6d0f71a73b75b9f15a05b3900811484d903e422c85f6
// 0xbedb226c3ba5e9214449d29319c3fea242e954e2f6c42c5dac56c300b61f4538
// 0x476f262f24f07c8c97354719605ac3137e341e9ba7dc63e9dbd342b2badf62d3
// 0x901513d973e19b594f3501460999b539e957f300fda939ac06df689590f6d206
// 0xaa30f5781425abb46471b997683171941b157cac093a81ad805903cb0d9fc946
// 0x7289736b6034fab8f4a0adb7c00281fbbbfe1c4b700d6c653c2bf77f71ea0dc6
// 0xf86abdee0b74ccb7c7d2e8db60a746475b4a94b7e4e12f4824192dc7031f3118
// 0xbce938c75d27abcb5774e84561808db4d56eb3c260c25dfcc9325b8be4b4bbf1
// 0x304c97d0fde7d8d40c45ed88964a121f2cf88b47eaee7e2f3884389b3ccb6a5d
// 0x4fd2a706afdc4a80c8f37217985ec9dfb11646c7d8c7b5656c03cdc42f9881d
// 0x34beebb6127e901faf99ac0ef87eebff71f8b26547d6cc8695d55bdeda8bde11
// 0x6713c45185cdbd3be7a22b3b0a59b071d9d9a30f97cc44886b7798d5ffa5cf20
// 0xcb739dd41e040ac96b849e1c5beddd3599ebc511cac1e1a605c5eedd6277a779
// 0x3e4c585eb0be545700305e26095d1a58bdafd2225bebcd49d3ba3c830ef2755e
// 0xc596d2eaeb9fba6cd6f1618dd62f0154a1599fffc1d5ccc7336adab2c5528e9
// 0xe5e09f9b2fd1df98e3b776285af5c278869d4d7955c2f6a8ea42dc61ea9b7995
// 0xdcd56b6f8a7b4f52516b93e6e030f139c7ff6269ea1e4ad9bc5e37b8f9cda0ba
// 0xd6cd761e99c2b63275dbd482cbf21b15b79406854cd06480ee5810439d89212a
// 0xb3cfcbd4ff2a1e55ec8a2ef5cc6fdaae19c20c9c65fc8f590f7794cabd57651d
// 0x3c388c700a2b8ba2530cf7bf0a30184de95c8bc49d473a3a38c8f39a4a0bb10e
// 0xc0bead20feada8bef3e6f4a12e4f409d6e4d636e3ed880ed9ae6e2255667c8ec
// 0x3bf16e19b3ab853d0d64695745544b38cd679d0e220f6b9c012fb54cd8c92334
// 0xc8b262d5c7b931ac993b84a051343ec74a7071ef37a95e16365b9639a1be5d3
// 0x4e84f2cb2665af7b42cc82f3a49482a8de03570bb25157a0503ef9ac6638f154
// 0xdcde06d9c4e8d9d1d77af05494313fa13a07f7108be2b861715c3c430cd6b4f7
// 0xa79a09a8ae75fdf46959f6f1ee938d3441ace7092d17b4c09f0a6d3103b5cf2e
// 0xa545ecf99aaa8ebf247691b97239b0cd45706d8ceeb969412a3c036093c5ed05
// 0xb83e47a153e664bf0224988d758f80e9dc2a524def60588bad71b7f18a52506
// 0x3ae855a18daadf9a6c0508a57fb4ad5055064fdd38a80831cd6fd5ce2513d8f9
// 0xedc33dbb416269f33bf2508fcbd68bf5312c6f9f1680c0e4513c71432c696e6c
// 0xee484b274efdb836cea9b09b9039226ef6dcf21467cc8a77486930fe28a9e17b
// 0xa77d7692a1e7eb7e2f507bd1718bf1eba8be8d006476a72f290fece9250a94ac
// 0xdd1f1721f880be6de850124a3ce0fa58f00da03d8af0f034cc124d96750b2943
// 0x4bcc4c059f41dc7574bea57e7f73d512685316d45b67cac93fa3026f6047823a
// 0x83d595f3fd1602ce40205165f1b824b57abeb4f1590a8e7e5e1bc70bf2462642
// 0x2ef9526bba21f8a025033f78ed9cb863c2a51a5942d8d4989ae698608a9417ab
// 0x38c30f133cf236f77b8f4bb6ac2964a96d73f6f36171a3d1cd0af2364289c351
// 0xc330ae25cf43305970b1b949d32223265bc16fa92c0995d17ef3e65d4d2ed1cd
// 0x6e2193eb2db96c81d584654a020a043301cc1c05d01593ab1a40178237f95171
// 0x27e944c3d71802cef21ad75806fbc23642fecfc5a7ac25060cd1e6180573d774
// 0xebdb696564f0b5f2b7a52d4b264eb1e1f2b9aa8699631412affef61bb1970418
// 0x49b5135f2e4958295dd7a32a9303998b17a20c5181ee7f783368c3cb65b16440
// 0xed466b635a15b1952454bcca1655042822a8d21079f7050fa7f3d47b330e2e1f
// 0x907ee22127ec6390aad4c384088af9c0d1a0f4d28b9d56b5d263bd0537c6fcb8
// 0x5e4bc4b76494fcb1ac64cda971a82c8cedef51cfad1dcc4d4278ac8098c2233
// 0x1ca62a269be9b36453a861c91c746d99ba33283a4cd53b86885c69d7b86d0ad7
// 0xc781d5f8f50ac9e54365ec2e5759aef039e1f0fe2664d967b18e72273bf2fddc
// 0xebe2d4ba89a720bca07e6ad55a5ca6480dab0bd8e7296777e7523fc306bbb9c
// 0x94e823d5df07dc672239d25875bf41316188b44ef55d889d9954fa1aeaa91477
// 0xf9dbf6affac9440fcbcdea210fcfe686ea86558ab506fc47773537b8b219d85
// 0x7001dd959f9360c4bd290c214d4690a14fee61dbb28ff560fbb77c74b1916ce9
// 0x958df0f64c724fe8612e2d0a818ae51c405e83cf1cbca85e7fed1dd0faf42a7e
// 0xff965948782d036c52e566f02edfae0c3e8a03b23fc590cbf3817ecae12b22f7
// 0x64b42821b68267504c685075f2ad7de806705db211c5c9e6889c00f4afdf9e1c
// 0xdab910a6721f03860a31083ad804a8bbf0e32e53684f8d4aa6c8142a31e39c54
// 0xd9640a3dae9c9088e5084ccca697775b0452feb130a5840722e1f311887caf6c
// 0xf3a5ee3a5dc8987dd7fba78d0730c6c88903073f2958f2bb9715bf1f202ee59a
// 0xdfacd83f20c4fa135f6746df0b4188a2d004efd68e8ca29c9365e2e904c742ab
// 0xe95c7fbfeef16cabc5f8d2ab9414d86449b50b873b308512a5f20e621f0dedee
// 0xc8860bd22d017dba93a1d35baed7b94ae6c4fc4900b3f1dd42d9c3de61cfa1dd
// 0xe903bf373e2f837ac8158c549179359e7a69b1143bb675f469ef82be8e4281b9
// 0x7824f8ba266763668d2f78edbb1c1d7b02c1d1bd5d22951882646759fb26600d
// 0xe57822ee7c6f22f3ae6a880505b15b3a09f28fc01868cbf8fbe98889ea7e1100
// 0x792454dfb432902ee5dd1846e4e72f822472a6d19edb9547c7a2663feaeb4f7a
// 0xf83a5efad7c764cefefa4335cda94721a76acf44512699000eca85ad2a77e59a
// 0xe827480a766b86abd48b50c7ee303d6a4469e508c141e83e8c9a3e0fead4a1ef
// 0x766293f6f81211a1d72c5c2c1a13681eaf42c57b46aa1bd6c5a50933e3df3040
// 0x34b382c8e1b123f751784d25294c7e53bafcfcbdb39fc4bbe6c3fa512f9d3ae7
// 0xdefdf14cf33e673c9e6107799a7bc4dc8024f2175c839ceb5f548a2672887848
// 0x60f4ff8282fffae3b12f443792e3ec8269ffab0117e25674fec223a525a5e8ed
// 0x294f143480f3b6dd37231bf69105456c9ca72cd657d7140fb7c1a8673e9d4c50
// 0x28a20c44bf10ee3d116950432c508c22f20890226610f4d8779347c5da460b18
// 0x377e51c14e788f1e22e4274b4f032eb9c396feb0be5987669440c3e1042d7f8c
// 0x65a1c9a048440571beb1a5f2357bc59907b69cc63f420f35a39bc2c80bcc4abe
// 0x56f99859bad886ff4c07a91621e651e99e622a168cb1c51ae393b8ab3c92482f
// 0x5662c33d851e4a1fb39111249b1bcfb8f3e2dd53930e16105fcf947101a0c1c7
// 0x7275ad80a7f16bbb972e8ddfe1b14f8300dae130b0cbdc241783e7415482e644
// 0xbd69bd2277b47ecdcd80381d8503521f55d4cdbd8901531cf8a3c81f237ea337
// 0xe24bc393cfae6feb1d51758476b1844ba882cbeb9cfd9695229d93c5cda36c1d
// 0xc4a007d214196436ae97e0254d34a0db7cd0c0a06b245c0dd95d2a22449e39b
// 0x49b956274e32b814db5a2f7b4f5e361e8bb459a9b49e8c2b9c0878f8bc6cc03c
// 0x3eb69851f836ae63467167b2943d1fd82840af6932929312e4a2b426fc6f2166
// 0x7bee29d373d29ae44bc19a688bfad497df082fd583722eb1d2924926292fc84b
// 0x4a3c2bff41ae4a9f554ecaeb865e84e791949f63b8680b9414dffe7c1cdc9419
// 0x8f6d1aa83120fa06c853eac2880eebb2902007813d7085ef0665c2a3cf67e0f1
// 0xe06e67e37a879f9da58c2346a89868f3924f3e0cc3a6436919fcfb3143cf226c
// 0xbd00350662bbdf968ab38a64dd8a7a86031815858d5bb49cd3f5a6dab8713217
// 0x977f5ec57cf100e526e963677de6301df44e2fbfb5e561efb0ea4b0a82b2de76
// 0x7890343258ebfafa1fd53cc14cde3e133cb4e5ee8706e8c7a0735333ca660ebb
// 0x36e68e7532c1f378289aef2fe8748f8e2d023682733da62b191306ed0ecb3226
// 0x3ac2839d8ae6d0ce0e61c331f0c8aebf384f511a267eeee67adf1aef9e7eff27
// 0xbd860e9ef67ef7ddb26be9d39d72c5a81c89f5ab4fe89e63b3608193a9a3915c
// 0x9aedb2a7d5f3539ee7be410865432548c0fcc5593cfc65d9a6f3f3ae6dd3d1f1
// 0xb3c9319cf12d4a4f791fcbda94209e7404845424fc87304453019e83997cdf4b
// 0x5d8b02613b4b2ee53f204ccb20d2650612da352703ece949385d86a400975a3
// 0x1728994ef17453728e51edd0e7d8cee9e864d84e50fb2a065cebbbeb1b1873cf
// 0x464de5eeab0b1f6526b911e95d4f68bc3a0426f5dc075141df311e0ea0bef841
// 0xbec88ca124a8a52851bd99784df633b8575c534b5c276369080e2c7385c71ae7
// 0xfd98a9243d2093792e5628aa9f3540d0d21592a734fff4d31f0037ea4da8497b
// 0x40fcecf7d38bbbb3905bb9d05b3cb88eb6d2dd051283b830e86d010938f11e4b
// 0xc87bddd3230c93be80e574eaf8bbaabd09c844268e73ca8ed76c1bc6369b42cf
// 0xcc7f0b15ec48305fe69aa7e2a0bd2ae2594f8d9906322beb4a9a40cdd9c1dda
// 0x38d0f34f8544f3d876c3771a1e80a3e61bee5328dac85805e54babc4bc2151b4
// 0x697735a831db03feafc74aedada2ef4285b875bae583ae88464ed82e3b8cdba
// 0x2292345a090754cedca733725c5ae81b5a922b59a60a84edb27e446e1b9b67af
// 0x7708d6ea813c95d3416e024a3ef3ccd1b8d2cd178b28ad50d15a9679c14a861b
// 0x3a536daaf751de5d88815b174e853aa602087244958fc7ffadae8d8cbd3cba05
// 0x49ab961254693024e3a955801e0c864be829cc09fb982b2cc5a8cdec35ff20c0
// 0x56eb8ff89c97f540da2aaea6e508d3b92e777a71a871620d09f8e5d44bdab6ab
// 0xf23d2b43ea37430f870cb3a759d1d4ec20a1c9b856592200a0c843b02b469866
// 0x8610dfaae52b9f26f354af75d776a87a645f05a8fe8c4f69512888cfd96a27cd
// 0x10f75d4f184384e40eefea494ecddf3cc0785f182db145646499ac6b1951729c
// 0x76a74e113de4538c60e8c40343486be360bced00f0b611280dbbd25f10ec414b
// 0xe955a760d68257768576f34a36890a2092227a7beb7b0b9551f0e7a8265570f6
// 0xc06d863c9baf4946ce555d51f572c24f05c5da24e388c3626d19e902a810d029
// 0x41b02617bea9f956f103aea1c922aebaffdacaf7567ad9f86048c7ef33934c29
// 0x54fbf23d3f1d580bef6ddd5dc8869df05fdd770fdee09842fab04e6c29f8f8ae
// 0xbffb89fa4a905c933e94468e23ccaa457af235e8a53e86debeedd401d6451946
// 0xb67094b5b1fb3c06c685d7c99468a53d88f066c9b29a3a222c3a451ac8b1e43a
// 0xe543131fed2faa58aa6c3606cc1e812b86ab5171ec35804a369cd22bb90f7953
// 0x37725ad61341fc5e12bb409ad97eee21fd4a1bfe953e790be81e9fc377d1e79e
// 0x1aac38954a51cb74b281a0781b810dd61b7e8a753d59ae30e4ac3208ac1bb3b4
// 0x41288660fbbb8a11fb3805d659e24f244d4a954e3bead32576fa24f59b108db4
// 0xc5311f3d23d086ea86f5ee7f85247b40896e29a0e251b00b0e2385aa114d6506
// 0xac3640ddbb2416e94e77b4a819d6344be01d03a35a9447d0c0ed447856ee6cc1
// 0xb5027d4fd9426822f2e67f6ae6cbe79505be5e4c8e7076320736f26142d6d278
// 0x40cd0923fdac9f0ac89d5137f1185797906029252fc007346391949fea5270dd
// 0x8c4a7723a566b5fbccc968a057dccda4156124d7251961dfa6ac66611b576b5a
// 0x53b18dbe9c58bfc66e26212ca02d4a03a26d0a0a4ae1dd52e9d6df265bfecb35
// 0x41cc680d1b995ed3db8ed0cc64ba3374d47e0c169dc28b2047bc206809569a33
// 0x232b3d76b32dad267e905125f621fd4fed644742578f22599472b0abf9dc5f8a
// 0x52cb7e443ff78d62e275551c75eb96b163b98e92d040c3d9ba3cba300044ec69
// 0xab2ebb74d7485e023d1705cc4ba56b62ed26040c67cff4441c673256cb676e06
// 0xec4fab731e2301ef164c0b26fc8fd88667d126d254229941d8412f09db8034fa
// 0xb81d40a1311014e81455983c79c8aa5d6a9a0791fea31dab5b241d379799b27a
// 0x79d9c89227487ecd478bbdfab355bbd5e4272022392dadf96b531cd975fa4171
// 0xced950ab9522026ea3b433a03ec8c0ee99dbf33fc414abc347e4e171cd440f13
// 0x1eed11e0679a40cdbf9ea05ae8c21bfe59271dce8da6476411b32dcee4136e38
// 0x3a2e8210702b55d9ec68adfa8be09ff224414a7a073259a9dff7201202f0b549
// 0xb20e58aa6fb2c054510a4f0d81fe55a07804beb5872e48095ad1f59a47fb118e
// 0xa04c8273003675f735cd2cf4092d14297c06cff6f2749746ccfa8fd2ce177870
// 0x902ddc82f7196ec79380cd92b4d37eeddf9ae6aff28ad4c3981b786fbd3ec5ae
// 0x415a6890434d0207a587e549a4926f68da2228f643777517ef8319bf0b8b8182
// 0x71cfca10bfe2dfef6ffb78f9141a4cd42a75fff8628cfcccecf159631dfab34b
// 0xeaa32a1319d0be3135ac92be6ee5a8fafe223ae4b916743ea8890bb198a6f16
// 0x37c1a0ed6fe0590667b160c4cc66754ee433e6dcfe219e7a2b43bb1b8ef1cef5
// 0xa3cce06c19044e99f9e915a77ead80d40d2e7a65fab2dab9a9389a69ec73bea6
// 0xf87fe8aaabe4f5e48ecea91a81e006029fecd1ed2932c23cc149cf9af560ddd
// 0x5403ac326bc7f12ea6b832c2abbc253bd415039e5b13960e47b49a05c5276dc7
// 0xc65afe6679d4665a4ac8586739b6c37b08319cc09ded9b798f7a165f81e329f2
// 0xcc58e6528d01979e5dc5cedcb5c25907ddd5b56fe4353bda1b03669cad7496f8
// 0x4f4000c5bf12be66290cf0e46b8d1d7abfac7580a78821c600823974e7b3f1b5
// 0x5b1a98d9b5b3cab3008545b480b0f0363657f78a8b0662278304138c71e376b1
// 0x7edbc5451cb634ce3d5d2e3d1d22c0cbe6c3ecf145fdd75307f8ff3d4ec8245d
// 0x404dee235637760b132777cd511015d01e24887252f8495d1b4556fd4f3fd8ac
// 0xd429a89fbbaa6c5078f8989968c68abb0c22fbb6bcabfbcf2499e037e579efc8
// 0x4aa9a5f75644e7e2ea634ea1a4787dbfc3e5e20660f4bf89b77936495e5d7123
// 0xba9c33b6b09b9603f588719907ea12bb629837aa7fa4944e9143e8965c32d1c7
// 0x8fa3743b26079d11a924758620ed8a3603731cb18ce896ba156024dd28e1fb65
// 0x2983f724a31f99054240d64f914e36dd1dd929919d5ff565fefb4f2fd0aeee01
// 0xefd987e5df91cd1596e0f84b635918e26d89dcba3123267df316e732ad179e18
// 0x7e8162b090e1cb38fa2234bd54eb6774f3337e47e962cf7ea5ca7d9ce4122c0d
// 0x3c6cd6a9b8fcba7f35b6868c465921cdf6018ae5c69fade42d4f70448b04dc18
// 0x42398692d2e8e97f285ed30b6d0864f5414f27abfec355982d997585d4a8ecd1
// 0xe184356e6b16120951a0260014ede9eca9248ade80c115228b1a0a7d26208df4
// 0xcfb586959347eff4209717612e8a08fc71ef35e04c2447d5018800e6cb1b8039
// 0xb1701069e2b9fcffd3d26f5e14f7b519df8147449c12d02e9efb2b0e57c48ed2
// 0xeb91c97362df6efd466b899b760f301da89fee596f6dfbbc9580390739b6dbaf
// 0xf87f7a0bb8b2709c6d7d7ee9ac64b335b5c95b5637f020fec7cee5121be61eb1
// 0x7fcf39de89f2872db4a5f565b320f6ed760017b135518c1d5b1b3b833e78ee7c
// 0x827e19e46434890ee62c9ca826fc40183e06339f5edef71a533d6222bcfaecee
// 0x6000305cc8e9cde03aad4a8dbd8fcea29871b6d2776f26cd54ccb96ebcf95709
// 0x6a8311c0d773bc48dfe0025da18359ff2fcf82cb3303e58f40794f6de518de7f
// 0xbd7b4761c3c434bdaf11cceca7aa19f1a84f98778c7ebd0236129d1913b84515
// 0x5966735305e652d38c52968f860f6e49cace832a9cb9be3711bc86b0f7fcf090
// 0xca74c64bffae5524e192b82c48210a1054d1183a0d0aff541a237b2ae48f5d62
// 0x89f339cf34dd9f779a153d2c758db89614b2d1518c0f96063383621c455b95c8
// 0xab4a3a487e8a7bcc952a53d459e8135fc99834e22ad8163df9331ef49f81078d
// 0x1f5e4ba770e9c1be392496c0d13487725acbf228dec9e1209020fa1c3b1ec961
// 0x39a5ead96290dfb4b213d13dde73e7fabbdad1ed9d7db73947200c5ebdddbae
// 0xf770d1e2507afa8c3e639e6b583771cfa3f6044ac0ce2475892281508df3d163
// 0xd98837040e7f7174f2fb78eb934e5732fae2c89101cce5ed67295d3fa2fd8e11
// 0xcb9b80ef91b09c5af530def5238d7fe035f71f52238f8ebe4882bea5ef13db6f
// 0xa19f4a81484404b056374ecf8b7e217936bc49a7929a7a37f6658f5c579736a4
// 0xe92ae219f2fa7897250eec27133d6efa151d47f40925a3cad834ef909f26666
// 0xffd8848a888bb4f5f430e6a81c8df9da76badb582195ef8ebd6c07a1fe985d85
// 0xfe16b23143dfeb977939f6e94976fe642433e34af1f62132a5e657bf3d1da5f7
// 0x8f5f007da4bcf5f2e1b257d4f566db7bf372d0ecd635dbb41863f5e83e608600
// 0x5a6a64907f2b26af5c2e8b05487449289384508f9ac5215527a2b9aa462cb6c6
// 0xca21681a8e34db51ef5bf608f5a6b49669c684a185d2ca93bb67357e36f873a1
// 0x8a6deb4343947b82eb6721ce3251c1190ecd16d8be3cdcec7e18e829d9617a4
// 0x3d0ba18f6e4affe6d0dd683923c1f25d3438969760f69b3c6da3fc0cf1224fb6
// 0xbedbcfe91d7f4d4779aa90c8e537c02624a4e6d78496938643433c75bf123622
// 0x799eb40085b64a98dddfb1a734c5c9784a110b563ffbc841ca4ee6589eac80b1
// 0x8006cccaf2a439d2769ace60351443168894d07e178bd8f029b2d43d948f3aa3
// 0xd73b3bdfa21ffeb8f93bf9b4c854279a0d5afdf0bcfeab0208d19f5a7ca89f9
// 0x4bb29ccf96fb21a3b3986e727eae30c5a383171772853f2157389588a91171d0
// 0xdb8ffddd3fdaf11fcfc4dfeac0e802d5f8acc994f31fcc8f14385c72f76b98d0
// 0x574388118b01f18e6c9da1a9d39e896ea9a2b4fb94fedfa28d9136acab9cf9cf
// 0x185ddf4e32b4ba43ae193fe8b7b3c2951374c86a1bcf934c31e0e7a8533b7d0a
// 0x8232dfdd35ba65851e5d0e9278dc6a22f1836b2af80efb3f75195eeb51f7ff05
// 0x1f327212e4c68b288b1b3b07af0f38663ba5da06a223395aca6ceeb82adc1eaa
// 0xe8662c4de2e75dc17ee1783d084476c1f1a51e280f3d9d0d41719933fb40dc37
// 0x2da137c68aa64686547046954b4fd7195dfe6784677a2fef86574738bafb71d2
// 0x8a4055126f108c4329695e526f6b723496e22db2d1e6e01dd550b39ce10d9702
// 0x315e45b7ca466267c3f869704ebee246a17ff179a03008ae91333f44f7364b60
// 0xfe088dbe324f0673c8b2cb4361b4d0d1e327074b5def36fab622fca4294c4859
// 0x55fe1512c9dc179b939415e0755d218912daad9d20f42c30173252dc819af1de
// 0xff7d3d1bfcfb79bc5f58f756f8c372554b4cf722d28f95b12ca6d60c370f8db3
// 0x9e9055711090c5b180a83b4b8cfffa484f61aed3f404c3564f167b7cab2b7722
// 0x3df9f187df65e0db9b585fb11c4b25b8046ef8c2a9f108c350b8cc720d76e89d
// 0xc012a5175f18b4bfb410691a1aa7c41fec35e174661c365e060b91d740896b00
// 0xfb978677b9b35accab1310024f645b5b4552fce0d75bb45fc083bf0038830430
// 0xb7aee50d7d8d6ee699c21c9952d9f5d3cd9f42403dd6201b7f28ab8133f72664
// 0x692c8f7d081cf958c631d6cbe7df5265a2b2962ed7aa329e78027ce425e5ec98
// 0x8ab797e3fb0ceb58f129fe853c9d5f38c58babe7b44f8e96db2fa1dd64911de7
// 0x93e16874891789ee1fe08e89890dffbed20a63aaaab3c133812bde92a2b79626
// 0xeb77c3adcae15b9a3146c15dbcefe2bcb62d2bed0869ace8e143a3f0db6e9a1d
// 0x62f784155fb4e0263bfedc8f0e60350101f80d67f3642b58816bcff3220e69a2
// 0x709b66d0ff01777007af055c6a0f80ebe1a9136c2a2cbeb9447414ab3a8f8d51
// 0x7a8b539d4b90778635ebaa7c89ac78dad98850c649a3cd68ca9f120acf523e98
// 0xecaef4d4695a11d272377e0d90f26414f902a7ef35f6f64fe5f7ac362374c819
// 0x7d166d724d00707ed3e587e70233c4572b219604496d2432a02e00a31454275a
// 0xcd9bd7ea9f2da28ca4063625056a9e060e726db60a9b7c7adb384a6a81b9a81f
// 0xfac408d9a40c255633c99b2b448485e12bcecb086077ef65dddfd21a7c31fbd7
// 0x24ba6b0249ed3c7159e86d0bd843068e3b15dc2c91ea8fb7629a49d36519a661
// 0xd2d7b733a2121a9176ba1ee169748bbc0e02eda2ec0cb90d7577c6ccfe058b4d
// 0xc8b5aa54533b64da5c45152680d6cf6bc3b10e0fbfec9e1f62343786cb43152c
// 0xc30c53bb3f36c4fbaaff4aaee5daf9277789d83ef7bc455243a55b311a73408f
// 0x3caf806d8aa677215e98464a97dbd84b4f4ebafb8c4d951d8a2b16d1c02b9616
// 0x92530b2e74fbe5e7280384c5bfa0f0722e8f64532023e5d354fa09a4e5813ec6
// 0x5023c56e0601f83ecef8b91c79af13cbf248e63145a76729fbcd7d6f263d1698
// 0xca43ac6558cb5fe49c6be40c37264ad818951a43d970b984283ae6d652eff69c
// 0xbfbde2ce6625324812543be5f23bcdb15bd4e82e3c49700e7e6393264c477846
// 0x7cc390e1f451bcc6af05560dc904649ca747d0f28a24bf75600162de71fc527e
// 0xa18c80e3b93a86d370cfef49ce429bd51b91bbe680420133c74ed7ec84e2f92e